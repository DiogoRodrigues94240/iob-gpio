   // GPIO
   input [15:0] gpio_sw,
   output [7:0] gpio_sseg_ca,
   output [3:0] gpio_sseg_an,
